module ioQueue #(
    // parameter
)(
    clk, rst,

    // Reqs
    reqValid,
    reqAddr,
    reqID,
    
    // Output bus
    rspValid,
    rspID
);



endmodule