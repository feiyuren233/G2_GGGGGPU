module name #(
    parameter FIFO_DEPTH = 16
)(
    clk, rstn

    // Req side
);
    
endmodule